* C:\Users\shree\eSim-Workspace\PN_Generation_ASHWINI\PN_Generation_ASHWINI.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 01/29/24 16:03:16

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ ? dff_sky		
U5  Net-_U1-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U5-Pad4_ ? dff_sky		
U6  Net-_U5-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U6-Pad4_ ? dff_sky		
U7  Net-_U6-Pad4_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U7-Pad4_ ? dff_sky		
U8  Net-_U1-Pad4_ Net-_U5-Pad4_ Net-_U6-Pad4_ Net-_U7-Pad4_ D1 D2 D3 D4 dac_bridge_4		
v2  clk GND pulse		
v1  rst GND pulse		
U12  D1 plot_v1		
U11  D2 plot_v1		
U10  D4 plot_v1		
U13  D3 plot_v1		
U9  Net-_U7-Pad4_ Net-_U5-Pad4_ Net-_U1-Pad1_ xor_sky		
U2  rst plot_v1		
U3  clk plot_v1		
scmode1  SKY130mode		
U4  rst clk Net-_U1-Pad3_ Net-_U1-Pad2_ adc_bridge_2		
U14  Net-_U1-Pad1_ xor_o dac_bridge_1		
U15  xor_o plot_v1		

.end
